//module reg_file(input LD_REG,
//input logic[2:0] DR,
//input[2:0] In_SR1,
//input[2:0] In_SR2,
//ouput
//
//)